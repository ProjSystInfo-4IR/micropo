
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity lc is
	Port (
			OPin : STD_LOGIC_VECTOR(4 downto 0);
			OPout : STD_LOGIC_VECTOR(4 downto 0);
			
		);
end lc;

architecture Behavioral of lc is

begin


end Behavioral;

