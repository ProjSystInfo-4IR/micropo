
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--use IEEE.NUMERIC_STD.ALL;

-- Uncomment the following library declaration if instantiating
-- any Xilinx primitives in this code.
--library UNISIM;
--use UNISIM.VComponents.all;

entity lc_mem is
	Port (
			OPin : in STD_LOGIC_VECTOR(3 downto 0);
			OPout : out STD_LOGIC
			
		);
end lc_mem;

architecture Behavioral of lc_mem is

begin


end Behavioral;

